//==============================================================================
//  Filename    : Read-Write Memory for instructions                                          
//  Designer    : Romain DUCHADEAU
//  Description : memory for instructions
//==============================================================================

