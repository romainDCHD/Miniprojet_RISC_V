library verilog;
use verilog.vl_types.all;
entity bench_control_logic is
end bench_control_logic;
